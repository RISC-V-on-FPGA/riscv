module uart_interface (
    ports
);
    
endmodule