`include "common.sv"

module decode_stage (
    input rst,
    input clk,
    input instruction_type instruction, // From program_memory
    input 
);
    
endmodule